module;
endmodule

module();
endmodule

module /**/ //
(/**/ //

) //
;
endmodule