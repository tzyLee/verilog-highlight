module _testbed_01$;
endmodule

module/**/test();
endmodule

module/**/ //
/**/ module_name
//
(/**/ //

) //
;
endmodule

module complex_ports ({c, d}, .e(f));
endmodule

module renamed_concat (.a({b, c}), f, .g(h[1]));
endmodule