module _testbed_01$;
endmodule

module/**/test();
endmodule

module/**/ //
/**/ module_name
//
(/**/ //

) //
;
endmodule